`timescale 1ns / 1ps    //Устанавливаем единицы времени: 1 нс, точность 1 пс
module jk_trigger_tb;
reg j;                  //описываем переменные
reg k;
reg clk;
wire q;
//далее необходимо подключить переменные
jk_trigger DUT(         //создаем экземпляр модуля 
    .j(j),
    .k(k),
    .clk(clk),
    .q(q));
//Далее настраиваем тактовый сигнал
always #5 clk = ~clk;   //создаем тактовый сигнал
//Теперь сам тест. Что и когда подавать на входы
//Начальные значения в блоке initial
initial 
begin
    clk = 0;
    j = 0;
    k = 0;
    #15;          //ожидание пары тактов

    //Теперь настройка j и k, их изменение увидим на следующем такте clk
    #10 j = 0; k = 0;   //хранение
    #10 j = 0; k = 1;   //сброс 
    #10 j = 1; k = 0;   //установка 
    #10 j = 0; k = 0;   //хранение 1
    #10 j = 1; k = 1;   //инверсия в 0
    #10 j = 1; k = 1;   //инверсия в 1
    #10 j = 1; k = 1;   //инверсия в 0

    #20 $display("Test complete");
    $finish;            //завершаем симуляцию
end
endmodule


