library verilog;
use verilog.vl_types.all;
entity t_trigger_tb is
end t_trigger_tb;
