library verilog;
use verilog.vl_types.all;
entity tb_gray_to_unary is
end tb_gray_to_unary;
