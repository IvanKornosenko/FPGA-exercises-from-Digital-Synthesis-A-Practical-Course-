module dec_6_64 (
    input [5:0] in,
    input en,
    output [63:0] out);

    assign out = en ? (1 << in) : 64'd0;  //Если en = 1, тогда у нас происходит сдвиг 1 на число in влево, иначе все 64 бита равны 0.
endmodule
/*Суть в том, что [5:0] это 6-и битный вход. В нем мы можем получить число от 0 до 63 в dec формате. 
  Для примера мы имеем 000111 на входе, это 7 в dec. Декодер делает сдвиг единицы на 7 цифр влево. 
  Мы получаем 0000000000000000000000000000000000000000000000000000000010000000. 
  Таким образом декодер активирует 7-ю шину из 64-х.        
  Нам это необходимо, так как иногда придется отключать и подключать разные устройства через такую вот шину. */
