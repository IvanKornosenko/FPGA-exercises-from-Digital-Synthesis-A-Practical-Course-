library verilog;
use verilog.vl_types.all;
entity jk_trigger_tb is
end jk_trigger_tb;
